module duck_hunt();

endmodule;
